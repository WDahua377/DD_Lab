module add6(a, b, sum, ov);

    input [5:0] a, b;
    output [6:0] sum;

    assign sum = a + b;

endmodule